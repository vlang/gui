module gui

pub const menu_separator_id = '__separator__'
pub const menu_subtitle_id = '__subtitle__'

// MenuItemCfg configures a menu-item.  Menu items are containers and are not limited
// to text. There are three types of menu items.
//
// - separator, if the separator field is true, a horizontal line separating menu items is rendered.
// - custom view, if a custom_view is supplied, it is rendered.
// - text only, for convenience, a text field is available for the typical text only menu items.
//
// If all three types are specified only one is rendered. The priority is separator, custom view, text only.
// Custom and text only menus can have a submenu.
//
// The optional action callback can be used to process menu clicks. There is also a catch-all
// action callback in [MenubarCfg](#MenubarCfg) that is called afterwards.
//
// It should go without saying, but menu-item id's need to be unique within a menubar config.
// This is necessary so callbacks can identify which menu-item was clicked. It also is how
// the menubar determines which menu items are selected/highlighted.
@[heap]
pub struct MenuItemCfg {
	color_select Color     = gui_theme.menubar_style.color_select
	text_style   TextStyle = gui_theme.menubar_style.text_style
	sizing       Sizing
	radius       f32 = gui_theme.menubar_style.radius_menu_item
	spacing      f32 = gui_theme.menubar_style.spacing_submenu
	disabled     bool
	selected     bool
pub:
	id          string @[required]
	text        string  = 'empty'
	padding     Padding = gui_theme.menubar_style.padding_menu_item
	action      fn (&MenuItemCfg, mut Event, mut Window) = unsafe { nil }
	submenu     []MenuItemCfg
	custom_view ?View
	separator   bool
}

fn menu_item(menubar_cfg MenubarCfg, item_cfg MenuItemCfg) View {
	return match item_cfg.separator {
		true {
			column(
				name:    'menu_item separator'
				id:      item_cfg.id
				height:  item_cfg.text_style.size / 2
				fill:    true
				sizing:  fill_fit
				padding: padding_none
				v_align: .middle
				content: [
					rectangle(
						height: 1
						color:  gui_theme.color_active
						sizing: fill_fit
					),
				]
			)
		}
		else {
			mut content := []View{cap: 1}
			unsafe { content.flags.set(.noslices) }
			if item_cfg.custom_view != none {
				content << item_cfg.custom_view
			} else {
				content << text(
					text:       item_cfg.text
					text_style: item_cfg.text_style
					mode:       .wrap
				)
			}
			column(
				name:     'menu_item'
				id:       item_cfg.id
				disabled: item_cfg.disabled
				color:    if item_cfg.selected {
					item_cfg.color_select
				} else {
					color_transparent
				}
				fill:     item_cfg.selected
				padding:  item_cfg.padding
				radius:   item_cfg.radius
				sizing:   item_cfg.sizing
				on_click: menubar_cfg.menu_item_click(item_cfg)
				spacing:  item_cfg.spacing
				on_hover: menubar_cfg.on_hover_item
				content:  content
			)
		}
	}
}

// menu_item_text is a convenience function for creating a simple text menu item
pub fn menu_item_text(id string, text string) MenuItemCfg {
	if id.len == 0 {
		panic("empty menu id's are invalid")
	}
	return MenuItemCfg{
		id:   id
		text: text
	}
}

// menu_separator is a convenience function for creating a menu separator
pub fn menu_separator() MenuItemCfg {
	return MenuItemCfg{
		id:        menu_separator_id
		separator: true
	}
}

// menu_subtitle subtitles
pub fn menu_subtitle(text string) MenuItemCfg {
	return MenuItemCfg{
		id:       menu_subtitle_id
		text:     text
		disabled: true
	}
}

// menu_submenu is a convenience function for creating a menu with an
// arrow symbol indicating a submenu
pub fn menu_submenu(id string, txt string, submenu []MenuItemCfg) MenuItemCfg {
	return MenuItemCfg{
		id:          id
		submenu:     submenu
		custom_view: row(
			padding: padding_none
			sizing:  fill_fit
			spacing: theme().spacing_large
			content: [
				text(text: txt, text_style: gui_theme.menubar_style.text_style),
				row(
					name:    'menu_submenu'
					h_align: .end
					sizing:  fill_fit
					padding: padding_none
					content: [
						text(
							text:       '›'
							text_style: gui_theme.menubar_style.text_style
						),
					]
				),
			]
		)
	}
}

// menu_item_click for such a short method, there is alot going on here in terms
// of state management, thus the many comments.
fn (cfg MenubarCfg) menu_item_click(item_cfg MenuItemCfg) fn (&Layout, mut Event, mut Window) {
	return fn [cfg, item_cfg] (_ &Layout, mut e Event, mut w Window) {
		// setting the focus to the menubar enables mouse hover highlighting of menu items.
		// see on_hover_item
		w.set_id_focus(cfg.id_focus)
		// Highlight the menu item
		w.view_state.menu_state[cfg.id_focus] = item_cfg.id
		// Menu item action handler
		if item_cfg.action != unsafe { nil } {
			item_cfg.action(item_cfg, mut e, mut w)
		}
		// Common menubar action handler
		cfg.action(item_cfg.id, mut e, mut w)
		// if this is simple menu-item (no submenu) then clicking it
		// also closes the menu and removes focus.
		if item_cfg.submenu.len == 0 {
			w.set_id_focus(0)
			w.view_state.menu_state[cfg.id_focus] = ''
		}
	}
}

fn (cfg &MenubarCfg) on_hover_item(mut layout Layout, mut _ Event, mut w Window) {
	// Mouse hover logic is covered here. Once the **menubar** gains focus,
	// mouse-overs can change the selected menu-item. Note: Selection
	// indicates highlighting, not focus. This is key to understanding menus.
	if layout.shape.id.len == 0 || layout.shape.disabled || !w.is_focus(cfg.id_focus) {
		return
	}
	w.view_state.menu_state[cfg.id_focus] = layout.shape.id
}
