module gui

// Based on Nic Barter's video of how Clay's UI algorithm works.
// https://www.youtube.com/watch?v=by9lQvpvMIc&t=1272s
//
import arrays
import gg

// layout_do executes a pipeline of functions to layout
// and position the Shapes of a ShapeTree
fn layout_do(mut layout ShapeTree, window Window) {
	layout_widths(mut layout)
	layout_flex_widths(mut layout)
	layout_wrap_text(mut layout, window.ui)
	layout_heights(mut layout)
	layout_flex_heights(mut layout)
	layout_positions(mut layout, 0, 0)

	width, height := window.window_size()
	layout_clipping_bounds(mut layout, width: width, height: height)
}

// layout_widths arranges a node's children Shapes horizontally. Only container
// nodes with a shape direction are arranged.
fn layout_widths(mut node ShapeTree) {
	for mut child in node.children {
		layout_widths(mut child)
		if node.shape.sizing.width != .fixed {
			match node.shape.direction {
				.left_to_right { node.shape.width += child.shape.width }
				.top_to_bottom { node.shape.width = f32_max(node.shape.width, child.shape.width) }
				.none {}
			}
			node.shape.width += node.shape.padding.left + node.shape.padding.right
			if node.shape.direction == .left_to_right {
				node.shape.width += node.shape.spacing * (node.children.len - 1)
			}
		}
	}
}

// layout_heights arranges a node's children Shapes vertically. Only container
// Shapes with a direction are arranged.
fn layout_heights(mut node ShapeTree) {
	for mut child in node.children {
		layout_heights(mut child)
		if node.shape.sizing.height != .fixed {
			match node.shape.direction {
				.top_to_bottom { node.shape.height += child.shape.height }
				.left_to_right { node.shape.height = f32_max(node.shape.height, child.shape.height) }
				.none {}
			}
			node.shape.height += node.shape.padding.top + node.shape.padding.bottom
			if node.shape.direction == .top_to_bottom {
				node.shape.height += node.shape.spacing * (node.children.len - 1)
			}
		}
	}
}

// layout_flex_widths manages the growing and shrinking of Shapes horizontally to satisfy
// a layout constraint
fn layout_flex_widths(mut node ShapeTree) {
	clamp := 100 // avoid infinite loop
	mut remaining_width := node.shape.width - node.shape.padding.left - node.shape.padding.right

	if node.shape.direction == .left_to_right {
		for mut child in node.children {
			remaining_width -= child.shape.width
		}
		// fence post spacing
		remaining_width -= (node.children.len - 1) * node.shape.spacing

		// Grow child elements
		idx := arrays.index_of_first(node.children, fn (_ int, n ShapeTree) bool {
			return n.shape.sizing.width == .flex
		})
		if idx < 0 {
			return
		}
		length := node.children.filter(it.shape.sizing.width == .flex).len

		// divide up the remaining flex widths by first growing
		// all the all the flex shapes to the same size (if possible)
		// and then distributing the remaining width to evenly.
		for i := 0; remaining_width > 0.1 && i < clamp; i++ {
			mut smallest := node.children[idx].shape.width
			mut second_smallest := f32(1000 * 1000)
			mut width_to_add := remaining_width

			for child in node.children {
				if child.shape.sizing.width == .flex {
					if child.shape.width < smallest {
						second_smallest = smallest
						smallest = child.shape.width
					}
					if child.shape.width > smallest {
						second_smallest = f32_min(second_smallest, child.shape.width)
						width_to_add = second_smallest - smallest
					}
				}
			}

			width_to_add = f32_min(width_to_add, remaining_width / length)

			for mut child in node.children {
				if child.shape.sizing.width == .flex {
					if child.shape.width == smallest {
						child.shape.width += width_to_add
						remaining_width -= width_to_add
					}
				}
			}
		}

		// Shrink if needed
		mut excluded := []string{}
		for i := 0; remaining_width < -0.1 && i < clamp; i++ {
			shrinkable := node.children.filter(it.shape.uid !in excluded)

			if shrinkable.len == 0 {
				return
			}

			mut largest := shrinkable[0].shape.width
			mut second_largest := f32(0)
			mut width_to_add := remaining_width

			for child in shrinkable {
				if child.shape.width > largest {
					second_largest = largest
					largest = child.shape.width
				}
				if child.shape.width < largest {
					second_largest = f32_max(second_largest, child.shape.width)
					width_to_add = second_largest - largest
				}
			}

			width_to_add = f32_max(width_to_add, remaining_width / shrinkable.len)

			for mut child in node.children {
				if child.shape.sizing.width == .flex {
					previous_width := child.shape.width
					if child.shape.width == largest {
						child.shape.width += width_to_add
						if child.shape.width <= child.shape.min_width {
							child.shape.width = child.shape.min_width
							excluded << child.shape.uid
						}
						remaining_width -= (child.shape.width - previous_width)
					}
				}
			}
		}
	} else if node.shape.direction == .top_to_bottom {
		for mut child in node.children {
			if child.shape.sizing.width == .flex {
				child.shape.width += (remaining_width - child.shape.width)
			}
		}
	}

	for mut child in node.children {
		layout_flex_widths(mut child)
	}
}

// layout_flex_heights manages the growing and shrinking of Shapes vertically to satisfy
// a layout constraint
fn layout_flex_heights(mut node ShapeTree) {
	mut remaining_height := node.shape.height - node.shape.padding.top - node.shape.padding.bottom

	if node.shape.direction == .top_to_bottom {
		for mut child in node.children {
			layout_flex_heights(mut child)
			remaining_height -= child.shape.height
		}

		// fence post spacing
		remaining_height -= (node.children.len - 1) * node.shape.spacing

		// Grow child elements
		idx := arrays.index_of_first(node.children, fn (_ int, n ShapeTree) bool {
			return n.shape.sizing.height == .flex
		})
		if idx < 0 {
			return
		}
		clamp := 100 // avoid infinite loop
		length := node.children.filter(it.shape.sizing.height == .flex).len

		// divide up the remaining flex hieghts by first growing
		// all the all the flex shape to the same size (if possible)
		// and then distributing the remaining height to evenly to
		// each
		for i := 0; remaining_height > 0.1 && i < clamp; i++ {
			mut smallest := node.children[idx].shape.height
			mut second_smallest := f32(1000 * 1000)
			mut height_to_add := remaining_height

			for child in node.children {
				if child.shape.sizing.height == .flex {
					if child.shape.height < smallest {
						second_smallest = smallest
						smallest = child.shape.height
					}
					if child.shape.height > smallest {
						second_smallest = f32_min(second_smallest, child.shape.height)
						height_to_add = second_smallest - smallest
					}
				}
			}

			height_to_add = f32_min(height_to_add, remaining_height / length)

			for mut child in node.children {
				if child.shape.sizing.height == .flex {
					if child.shape.height == smallest {
						child.shape.height += height_to_add
						remaining_height -= height_to_add
					}
				}
			}
		}
	} else if node.shape.direction == .left_to_right {
		for mut child in node.children {
			if child.shape.sizing.height == .flex {
				child.shape.height += (remaining_height - child.shape.height)
			}
		}
	}

	for mut child in node.children {
		layout_flex_heights(mut child)
	}
}

// layout_wrap_text is called after all widths in a ShapeTree are determined.
// Wrapping text can change the height of an Shape, which is why this is called
// before computing Shape heights
fn layout_wrap_text(mut node ShapeTree, ctx gg.Context) {
	text_wrap(mut node.shape, ctx)
	for mut child in node.children {
		layout_wrap_text(mut child, ctx)
	}
}

// layout_positions sets the positions of all Shapes in the ShapeTreee.
// It also handles alignment (soon)
fn layout_positions(mut node ShapeTree, offset_x f32, offset_y f32) {
	node.shape.x += offset_x
	node.shape.y += offset_y

	spacing := node.shape.spacing
	direction := node.shape.direction

	mut x := node.shape.x + node.shape.padding.left
	mut y := node.shape.y + node.shape.padding.top

	for mut child in node.children {
		layout_positions(mut child, x, y)
		match direction {
			.left_to_right { x += child.shape.width + spacing }
			.top_to_bottom { y += child.shape.height + spacing }
			.none {}
		}
	}
}

// layout_clipping_bounds ensures that Shapes do not draw outside the parent
// Shape container.
fn layout_clipping_bounds(mut node ShapeTree, bounds gg.Rect) {
	nb := match node.shape.type == .container {
		true {
			bw := bounds.x + bounds.width
			nw := node.shape.x + node.shape.width
			bh := bounds.y + bounds.height
			nh := node.shape.y + node.shape.height

			gg.Rect{
				x:      if bw < nw { bounds.x } else { node.shape.x }
				y:      if bh < nh { bounds.y } else { node.shape.y }
				width:  if bw < nw { bounds.width } else { node.shape.width }
				height: if bh < nh { bounds.height } else { node.shape.height }
			}
		}
		else {
			bounds
		}
	}
	for mut child in node.children {
		child.shape.bounds = nb
		layout_clipping_bounds(mut child, nb)
	}
}
