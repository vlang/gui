module titlebar

pub fn set_dark_mode(dark bool) {}
