@[has_globals]
module gui

__global gui_theme = theme_dark

pub const version = '0.1.0'
pub const app_title = 'GUI'
