module titlebar

pub fn set_mode(dark bool) {}
