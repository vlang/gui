module gui

pub const version = '0.1.0'
pub const app_title = 'GUI'
