module gui

import gg

pub struct MouseEvent {
	mouse_x      f32
	mouse_y      f32
	mouse_button gg.MouseButton
}
