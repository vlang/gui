module gui

import os

pub const icon_font_file = os.join_path(os.data_dir(), 'gui_feathericon.ttf')

fn install_icon_font() {
	icon_font := $embed_file('assets/feathericon.ttf')
	if !os.exists(icon_font_file) {
		os.write_file(icon_font_file, icon_font.to_string()) or {}
	}
}

pub const icons_map = {
	'icon_arrow_down':              '\uf100'
	'icon_arrow_left':              '\uf101'
	'icon_arrow_right':             '\uf102'
	'icon_arrow_up':                '\uf103'
	'icon_artboard':                '\uf104'
	'icon_bar':                     '\uf105'
	'icon_bar_chart':               '\uf106'
	'icon_beer':                    '\uf107'
	'icon_bell':                    '\uf108'
	'icon_book':                    '\uf109'
	'icon_browser':                 '\uf10b'
	'icon_brush':                   '\uf10c'
	'icon_bug':                     '\uf10d'
	'icon_building':                '\uf10e'
	'icon_calendar':                '\uf10f'
	'icon_camera':                  '\uf110'
	'icon_check':                   '\uf111'
	'icon_clock':                   '\uf113'
	'icon_close':                   '\uf114'
	'icon_cloud':                   '\uf115'
	'icon_cocktail':                '\uf116'
	'icon_code':                    '\uf117'
	'icon_columns':                 '\uf118'
	'icon_comment':                 '\uf119'
	'icon_commenting':              '\uf11a'
	'icon_comments':                '\uf11b'
	'icon_desktop':                 '\uf11d'
	'icon_diamond':                 '\uf11e'
	'icon_disabled':                '\uf11f'
	'icon_download':                '\uf120'
	'icon_drop_down':               '\uf121'
	'icon_drop_left':               '\uf122'
	'icon_drop_right':              '\uf123'
	'icon_drop_up':                 '\uf124'
	'icon_elipsis_h':               '\uf125'
	'icon_elipsis_v':               '\uf126'
	'icon_eye':                     '\uf127'
	'icon_feed':                    '\uf128'
	'icon_flag':                    '\uf129'
	'icon_folder':                  '\uf12a'
	'icon_fork':                    '\uf12b'
	'icon_globe':                   '\uf12c'
	'icon_hash':                    '\uf12d'
	'icon_heart':                   '\uf12e'
	'icon_home':                    '\uf12f'
	'icon_info':                    '\uf130'
	'icon_key':                     '\uf131'
	'icon_keyboard':                '\uf132'
	'icon_laptop':                  '\uf133'
	'icon_layout':                  '\uf134'
	'icon_line_chart':              '\uf135'
	'icon_link':                    '\uf136'
	'icon_link_external':           '\uf137'
	'icon_location':                '\uf138'
	'icon_lock':                    '\uf139'
	'icon_login':                   '\uf13a'
	'icon_logout':                  '\uf13b'
	'icon_mail':                    '\uf13c'
	'icon_medal':                   '\uf13d'
	'icon_megaphone':               '\uf13e'
	'icon_minus':                   '\uf140'
	'icon_mobile':                  '\uf141'
	'icon_mouse':                   '\uf142'
	'icon_pencil':                  '\uf144'
	'icon_phone':                   '\uf145'
	'icon_pie_chart':               '\uf146'
	'icon_pizza':                   '\uf147'
	'icon_plus':                    '\uf148'
	'icon_prototype':               '\uf149'
	'icon_question':                '\uf14a'
	'icon_quote_left':              '\uf14b'
	'icon_quote_right':             '\uf14c'
	'icon_rocket':                  '\uf14d'
	'icon_search':                  '\uf14e'
	'icon_share':                   '\uf14f'
	'icon_sitemap':                 '\uf150'
	'icon_star':                    '\uf151'
	'icon_tablet':                  '\uf152'
	'icon_tag':                     '\uf153'
	'icon_terminal':                '\uf154'
	'icon_ticket':                  '\uf155'
	'icon_tiled':                   '\uf156'
	'icon_trash':                   '\uf157'
	'icon_trophy':                  '\uf158'
	'icon_upload':                  '\uf159'
	'icon_user':                    '\uf15a'
	'icon_user_plus':               '\uf15b'
	'icon_users':                   '\uf15c'
	'icon_vector':                  '\uf15d'
	'icon_video':                   '\uf15e'
	'icon_warning':                 '\uf15f'
	'icon_wine_glass':              '\uf161'
	'icon_wrench':                  '\uf162'
	'icon_birthday_cake':           '\uf163'
	'icon_mention':                 '\uf164'
	'icon_palette':                 '\uf165'
	'icon_coffee':                  '\uf166'
	'icon_heart_o':                 '\uf167'
	'icon_star_o':                  '\uf168'
	'icon_unlock':                  '\uf169'
	'icon_search_minus':            '\uf16a'
	'icon_search_plus':             '\uf16b'
	'icon_user_minus':              '\uf16c'
	'icon_map':                     '\uf16d'
	'icon_export':                  '\uf16e'
	'icon_import':                  '\uf16f'
	'icon_bookmark':                '\uf170'
	'icon_print':                   '\uf171'
	'icon_shield':                  '\uf172'
	'icon_filter':                  '\uf173'
	'icon_feather':                 '\uf174'
	'icon_music':                   '\uf175'
	'icon_folder_open':             '\uf176'
	'icon_magic':                   '\uf177'
	'icon_paper_plane':             '\uf178'
	'icon_bold':                    '\uf179'
	'icon_italic':                  '\uf17a'
	'icon_text_size':               '\uf17b'
	'icon_list_bullet':             '\uf17c'
	'icon_list_order':              '\uf17d'
	'icon_list_task':               '\uf17e'
	'icon_edit':                    '\uf17f'
	'icon_backward':                '\uf180'
	'icon_compress':                '\uf181'
	'icon_eject':                   '\uf182'
	'icon_expand':                  '\uf183'
	'icon_fast_backward':           '\uf184'
	'icon_fast_forward':            '\uf185'
	'icon_forward':                 '\uf186'
	'icon_pause':                   '\uf187'
	'icon_play':                    '\uf188'
	'icon_random':                  '\uf189'
	'icon_stop':                    '\uf18b'
	'icon_layer':                   '\uf18c'
	'icon_headphone':               '\uf18e'
	'icon_plug':                    '\uf18f'
	'icon_usb':                     '\uf190'
	'icon_gamepad':                 '\uf191'
	'icon_loop':                    '\uf192'
	'icon_sync':                    '\uf194'
	'icon_align_center':            '\uf195'
	'icon_align_left':              '\uf196'
	'icon_align_right':             '\uf197'
	'icon_app_menu':                '\uf198'
	'icon_audio_player':            '\uf199'
	'icon_check_circle':            '\uf19a'
	'icon_check_circle_o':          '\uf19b'
	'icon_check_verified':          '\uf19c'
	'icon_cutlery':                 '\uf19d'
	'icon_delete_link':             '\uf19e'
	'icon_document':                '\uf19f'
	'icon_equalizer':               '\uf1a0'
	'icon_file_excel':              '\uf1a2'
	'icon_file_powerpoint':         '\uf1a3'
	'icon_file_word':               '\uf1a4'
	'icon_gear':                    '\uf1a5'
	'icon_insert_link':             '\uf1a6'
	'icon_kitchen_cooker':          '\uf1a7'
	'icon_money':                   '\uf1a8'
	'icon_picture':                 '\uf1a9'
	'icon_pot':                     '\uf1aa'
	'icon_speaker':                 '\uf1ab'
	'icon_table':                   '\uf1ac'
	'icon_timeline':                '\uf1ad'
	'icon_underline':               '\uf1ae'
	'icon_watch':                   '\uf1af'
	'icon_watch_alt':               '\uf1b0'
	'icon_file':                    '\uf1b1'
	'icon_file_audio':              '\uf1b2'
	'icon_file_image':              '\uf1b3'
	'icon_file_movie':              '\uf1b4'
	'icon_file_zip':                '\uf1b5'
	'icon_angry':                   '\uf1b6'
	'icon_cry':                     '\uf1b7'
	'icon_disappointed':            '\uf1b8'
	'icon_frowing':                 '\uf1b9'
	'icon_open_mouth':              '\uf1ba'
	'icon_rage':                    '\uf1bb'
	'icon_smile':                   '\uf1bc'
	'icon_smile_alt':               '\uf1bd'
	'icon_tired':                   '\uf1be'
	'icon_align_bottom':            '\uf1bf'
	'icon_align_top':               '\uf1c0'
	'icon_align_vertically':        '\uf1c1'
	'icon_crop':                    '\uf1c2'
	'icon_difference':              '\uf1c3'
	'icon_distribute_vertically':   '\uf1c5'
	'icon_eraser':                  '\uf1c6'
	'icon_intersect':               '\uf1c7'
	'icon_mask':                    '\uf1c8'
	'icon_scale':                   '\uf1c9'
	'icon_subtract':                '\uf1ca'
	'icon_text_align_center':       '\uf1cb'
	'icon_text_align_left':         '\uf1cc'
	'icon_text_align_right':        '\uf1cd'
	'icon_union':                   '\uf1ce'
	'icon_distribute_horizontally': '\uf1cf'
	'icon_step_backward':           '\uf1d0'
	'icon_step_forward':            '\uf1d1'
	'icon_comment_o':               '\uf1d2'
	'icon_codepen':                 '\uf1d3'
	'icon_facebook':                '\uf1d4'
	'icon_git':                     '\uf1d5'
	'icon_github':                  '\uf1d6'
	'icon_github_alt':              '\uf1d7'
	'icon_google':                  '\uf1d8'
	'icon_google_plus':             '\uf1d9'
	'icon_instagram':               '\uf1da'
	'icon_pinterest':               '\uf1db'
	'icon_pocket':                  '\uf1dc'
	'icon_twitter':                 '\uf1dd'
	'icon_wordpress':               '\uf1de'
	'icon_wordpress_alt':           '\uf1df'
	'icon_youtube':                 '\uf1e0'
	'icon_messanger':               '\uf1e1'
	'icon_activity':                '\uf1e2'
	'icon_bolt':                    '\uf1e3'
	'icon_picture_square':          '\uf1e4'
	'icon_text_align_justify':      '\uf1e5'
	'icon_add_cart':                '\uf1e6'
	'icon_cage':                    '\uf1e7'
	'icon_cart':                    '\uf1e8'
	'icon_credit_card':             '\uf1e9'
	'icon_gift':                    '\uf1ea'
	'icon_remove_cart':             '\uf1eb'
	'icon_shopping_bag':            '\uf1ec'
	'icon_truck':                   '\uf1ed'
	'icon_wallet':                  '\uf1ee'
	'icon_moon':                    '\uf1ef'
	'icon_sunny_o':                 '\uf1f0'
	'icon_sunrise':                 '\uf1f1'
	'icon_umbrella':                '\uf1f2'
	'icon_target':                  '\uf1f3'
	'icon_smile_plus':              '\uf1f5'
	'icon_smile_heart':             '\uf1f6'
	'icon_beginner':                '\uf1f7'
	'icon_train':                   '\uf1f8'
	'icon_donut':                   '\uf1f9'
	'icon_rice_cracker':            '\uf1fa'
	'icon_apron':                   '\uf1fb'
	'icon_octpus':                  '\uf1fc'
	'icon_squid':                   '\uf1fd'
	'icon_bus':                     '\uf1fe'
	'icon_car':                     '\uf1ff'
	'icon_notice_active':           '\uf200'
	'icon_notice_off':              '\uf201'
	'icon_notice_on':               '\uf202'
	'icon_notice_push':             '\uf203'
	'icon_taxi':                    '\uf204'
	'icon_vr':                      '\uf205'
	'icon_bread':                   '\uf206'
	'icon_frying_pan':              '\uf207'
	'icon_mitarashi_dango':         '\uf208'
	'icon_tumbler_glass':           '\uf209'
	'icon_yaki_dango':              '\uf20a'
}

pub const icon_arrow_down = '\uf100'
pub const icon_arrow_left = '\uf101'
pub const icon_arrow_right = '\uf102'
pub const icon_arrow_up = '\uf103'
pub const icon_artboard = '\uf104'
pub const icon_bar = '\uf105'
pub const icon_bar_chart = '\uf106'
pub const icon_beer = '\uf107'
pub const icon_bell = '\uf108'
pub const icon_book = '\uf109'
pub const icon_browser = '\uf10b'
pub const icon_brush = '\uf10c'
pub const icon_bug = '\uf10d'
pub const icon_building = '\uf10e'
pub const icon_calendar = '\uf10f'
pub const icon_camera = '\uf110'
pub const icon_check = '\uf111'
pub const icon_clock = '\uf113'
pub const icon_close = '\uf114'
pub const icon_cloud = '\uf115'
pub const icon_cocktail = '\uf116'
pub const icon_code = '\uf117'
pub const icon_columns = '\uf118'
pub const icon_comment = '\uf119'
pub const icon_commenting = '\uf11a'
pub const icon_comments = '\uf11b'
pub const icon_desktop = '\uf11d'
pub const icon_diamond = '\uf11e'
pub const icon_disabled = '\uf11f'
pub const icon_download = '\uf120'
pub const icon_drop_down = '\uf121'
pub const icon_drop_left = '\uf122'
pub const icon_drop_right = '\uf123'
pub const icon_drop_up = '\uf124'
pub const icon_elipsis_h = '\uf125'
pub const icon_elipsis_v = '\uf126'
pub const icon_eye = '\uf127'
pub const icon_feed = '\uf128'
pub const icon_flag = '\uf129'
pub const icon_folder = '\uf12a'
pub const icon_fork = '\uf12b'
pub const icon_globe = '\uf12c'
pub const icon_hash = '\uf12d'
pub const icon_heart = '\uf12e'
pub const icon_home = '\uf12f'
pub const icon_info = '\uf130'
pub const icon_key = '\uf131'
pub const icon_keyboard = '\uf132'
pub const icon_laptop = '\uf133'
pub const icon_layout = '\uf134'
pub const icon_line_chart = '\uf135'
pub const icon_link = '\uf136'
pub const icon_link_external = '\uf137'
pub const icon_location = '\uf138'
pub const icon_lock = '\uf139'
pub const icon_login = '\uf13a'
pub const icon_logout = '\uf13b'
pub const icon_mail = '\uf13c'
pub const icon_medal = '\uf13d'
pub const icon_megaphone = '\uf13e'
pub const icon_minus = '\uf140'
pub const icon_mobile = '\uf141'
pub const icon_mouse = '\uf142'
pub const icon_pencil = '\uf144'
pub const icon_phone = '\uf145'
pub const icon_pie_chart = '\uf146'
pub const icon_pizza = '\uf147'
pub const icon_plus = '\uf148'
pub const icon_prototype = '\uf149'
pub const icon_question = '\uf14a'
pub const icon_quote_left = '\uf14b'
pub const icon_quote_right = '\uf14c'
pub const icon_rocket = '\uf14d'
pub const icon_search = '\uf14e'
pub const icon_share = '\uf14f'
pub const icon_sitemap = '\uf150'
pub const icon_star = '\uf151'
pub const icon_tablet = '\uf152'
pub const icon_tag = '\uf153'
pub const icon_terminal = '\uf154'
pub const icon_ticket = '\uf155'
pub const icon_tiled = '\uf156'
pub const icon_trash = '\uf157'
pub const icon_trophy = '\uf158'
pub const icon_upload = '\uf159'
pub const icon_user = '\uf15a'
pub const icon_user_plus = '\uf15b'
pub const icon_users = '\uf15c'
pub const icon_vector = '\uf15d'
pub const icon_video = '\uf15e'
pub const icon_warning = '\uf15f'
pub const icon_wine_glass = '\uf161'
pub const icon_wrench = '\uf162'
pub const icon_birthday_cake = '\uf163'
pub const icon_mention = '\uf164'
pub const icon_palette = '\uf165'
pub const icon_coffee = '\uf166'
pub const icon_heart_o = '\uf167'
pub const icon_star_o = '\uf168'
pub const icon_unlock = '\uf169'
pub const icon_search_minus = '\uf16a'
pub const icon_search_plus = '\uf16b'
pub const icon_user_minus = '\uf16c'
pub const icon_map = '\uf16d'
pub const icon_export = '\uf16e'
pub const icon_import = '\uf16f'
pub const icon_bookmark = '\uf170'
pub const icon_print = '\uf171'
pub const icon_shield = '\uf172'
pub const icon_filter = '\uf173'
pub const icon_feather = '\uf174'
pub const icon_music = '\uf175'
pub const icon_folder_open = '\uf176'
pub const icon_magic = '\uf177'
pub const icon_paper_plane = '\uf178'
pub const icon_bold = '\uf179'
pub const icon_italic = '\uf17a'
pub const icon_text_size = '\uf17b'
pub const icon_list_bullet = '\uf17c'
pub const icon_list_order = '\uf17d'
pub const icon_list_task = '\uf17e'
pub const icon_edit = '\uf17f'
pub const icon_backward = '\uf180'
pub const icon_compress = '\uf181'
pub const icon_eject = '\uf182'
pub const icon_expand = '\uf183'
pub const icon_fast_backward = '\uf184'
pub const icon_fast_forward = '\uf185'
pub const icon_forward = '\uf186'
pub const icon_pause = '\uf187'
pub const icon_play = '\uf188'
pub const icon_random = '\uf189'
pub const icon_stop = '\uf18b'
pub const icon_layer = '\uf18c'
pub const icon_headphone = '\uf18e'
pub const icon_plug = '\uf18f'
pub const icon_usb = '\uf190'
pub const icon_gamepad = '\uf191'
pub const icon_loop = '\uf192'
pub const icon_sync = '\uf194'
pub const icon_align_center = '\uf195'
pub const icon_align_left = '\uf196'
pub const icon_align_right = '\uf197'
pub const icon_app_menu = '\uf198'
pub const icon_audio_player = '\uf199'
pub const icon_check_circle = '\uf19a'
pub const icon_check_circle_o = '\uf19b'
pub const icon_check_verified = '\uf19c'
pub const icon_cutlery = '\uf19d'
pub const icon_delete_link = '\uf19e'
pub const icon_document = '\uf19f'
pub const icon_equalizer = '\uf1a0'
pub const icon_file_excel = '\uf1a2'
pub const icon_file_powerpoint = '\uf1a3'
pub const icon_file_word = '\uf1a4'
pub const icon_gear = '\uf1a5'
pub const icon_insert_link = '\uf1a6'
pub const icon_kitchen_cooker = '\uf1a7'
pub const icon_money = '\uf1a8'
pub const icon_picture = '\uf1a9'
pub const icon_pot = '\uf1aa'
pub const icon_speaker = '\uf1ab'
pub const icon_table = '\uf1ac'
pub const icon_timeline = '\uf1ad'
pub const icon_underline = '\uf1ae'
pub const icon_watch = '\uf1af'
pub const icon_watch_alt = '\uf1b0'
pub const icon_file = '\uf1b1'
pub const icon_file_audio = '\uf1b2'
pub const icon_file_image = '\uf1b3'
pub const icon_file_movie = '\uf1b4'
pub const icon_file_zip = '\uf1b5'
pub const icon_angry = '\uf1b6'
pub const icon_cry = '\uf1b7'
pub const icon_disappointed = '\uf1b8'
pub const icon_frowing = '\uf1b9'
pub const icon_open_mouth = '\uf1ba'
pub const icon_rage = '\uf1bb'
pub const icon_smile = '\uf1bc'
pub const icon_smile_alt = '\uf1bd'
pub const icon_tired = '\uf1be'
pub const icon_align_bottom = '\uf1bf'
pub const icon_align_top = '\uf1c0'
pub const icon_align_vertically = '\uf1c1'
pub const icon_crop = '\uf1c2'
pub const icon_difference = '\uf1c3'
pub const icon_distribute_vertically = '\uf1c5'
pub const icon_eraser = '\uf1c6'
pub const icon_intersect = '\uf1c7'
pub const icon_mask = '\uf1c8'
pub const icon_scale = '\uf1c9'
pub const icon_subtract = '\uf1ca'
pub const icon_text_align_center = '\uf1cb'
pub const icon_text_align_left = '\uf1cc'
pub const icon_text_align_right = '\uf1cd'
pub const icon_union = '\uf1ce'
pub const icon_distribute_horizontally = '\uf1cf'
pub const icon_step_backward = '\uf1d0'
pub const icon_step_forward = '\uf1d1'
pub const icon_comment_o = '\uf1d2'
pub const icon_codepen = '\uf1d3'
pub const icon_facebook = '\uf1d4'
pub const icon_git = '\uf1d5'
pub const icon_github = '\uf1d6'
pub const icon_github_alt = '\uf1d7'
pub const icon_google = '\uf1d8'
pub const icon_google_plus = '\uf1d9'
pub const icon_instagram = '\uf1da'
pub const icon_pinterest = '\uf1db'
pub const icon_pocket = '\uf1dc'
pub const icon_twitter = '\uf1dd'
pub const icon_wordpress = '\uf1de'
pub const icon_wordpress_alt = '\uf1df'
pub const icon_youtube = '\uf1e0'
pub const icon_messanger = '\uf1e1'
pub const icon_activity = '\uf1e2'
pub const icon_bolt = '\uf1e3'
pub const icon_picture_square = '\uf1e4'
pub const icon_text_align_justify = '\uf1e5'
pub const icon_add_cart = '\uf1e6'
pub const icon_cage = '\uf1e7'
pub const icon_cart = '\uf1e8'
pub const icon_credit_card = '\uf1e9'
pub const icon_gift = '\uf1ea'
pub const icon_remove_cart = '\uf1eb'
pub const icon_shopping_bag = '\uf1ec'
pub const icon_truck = '\uf1ed'
pub const icon_wallet = '\uf1ee'
pub const icon_moon = '\uf1ef'
pub const icon_sunny_o = '\uf1f0'
pub const icon_sunrise = '\uf1f1'
pub const icon_umbrella = '\uf1f2'
pub const icon_target = '\uf1f3'
pub const icon_smile_plus = '\uf1f5'
pub const icon_smile_heart = '\uf1f6'
pub const icon_beginner = '\uf1f7'
pub const icon_train = '\uf1f8'
pub const icon_donut = '\uf1f9'
pub const icon_rice_cracker = '\uf1fa'
pub const icon_apron = '\uf1fb'
pub const icon_octpus = '\uf1fc'
pub const icon_squid = '\uf1fd'
pub const icon_bus = '\uf1fe'
pub const icon_car = '\uf1ff'
pub const icon_notice_active = '\uf200'
pub const icon_notice_off = '\uf201'
pub const icon_notice_on = '\uf202'
pub const icon_notice_push = '\uf203'
pub const icon_taxi = '\uf204'
pub const icon_vr = '\uf205'
pub const icon_bread = '\uf206'
pub const icon_frying_pan = '\uf207'
pub const icon_mitarashi_dango = '\uf208'
pub const icon_tumbler_glass = '\uf209'
pub const icon_yaki_dango = '\uf20a'
