module gui

const feather_icons = {
	'activity':           '\uE900'
	'airplay':            '\uE901'
	'alert-circle':       '\uE902'
	'alert-octagon':      '\uE903'
	'alert-triangle':     '\uE904'
	'align-center':       '\uE905'
	'align-justify':      '\uE906'
	'align-left':         '\uE907'
	'align-right':        '\uE908'
	'anchor':             '\uE909'
	'aperture':           '\uE90A'
	'archive':            '\uE90B'
	'arrow-down':         '\uE90C'
	'arrow-down-circle':  '\uE90D'
	'arrow-down-left':    '\uE90E'
	'arrow-down-right':   '\uE90F'
	'arrow-left':         '\uE910'
	'arrow-left-circle':  '\uE911'
	'arrow-right':        '\uE912'
	'arrow-right-circle': '\uE913'
	'arrow-up':           '\uE914'
	'arrow-up-circle':    '\uE915'
	'arrow-up-left':      '\uE916'
	'arrow-up-right':     '\uE917'
	'at-sign':            '\uE918'
	'award':              '\uE919'
	'bar-chart':          '\uE91A'
	'bar-chart-2':        '\uE91B'
	'battery':            '\uE91C'
	'battery-charging':   '\uE91D'
	'bell':               '\uE91E'
	'bell-off':           '\uE91F'
	'bluetooth':          '\uE920'
	'bold':               '\uE921'
	'book':               '\uE922'
	'book-open':          '\uE923'
	'bookmark':           '\uE924'
	'box':                '\uE925'
	'briefcase':          '\uE926'
	'calendar':           '\uE927'
	'camera':             '\uE928'
	'camera-off':         '\uE929'
	'cast':               '\uE92A'
	'check':              '\uE92B'
	'check-circle':       '\uE92C'
	'check-square':       '\uE92D'
	'chevron-down':       '\uE92E'
	'chevron-left':       '\uE92F'
	'chevron-right':      '\uE930'
	'chevron-up':         '\uE931'
	'chevrons-down':      '\uE932'
	'chevrons-left':      '\uE933'
	'chevrons-right':     '\uE934'
	'chevrons-up':        '\uE935'
	'chrome':             '\uE936'
	'circle':             '\uE937'
	'clipboard':          '\uE938'
	'clock':              '\uE939'
	'cloud':              '\uE93A'
	'cloud-drizzle':      '\uE93B'
	'cloud-lightning':    '\uE93C'
	'cloud-off':          '\uE93D'
	'cloud-rain':         '\uE93E'
	'cloud-snow':         '\uE93F'
	'code':               '\uE940'
	'codepen':            '\uE941'
	'codesandbox':        '\uE942'
	'coffee':             '\uE943'
	'columns':            '\uE944'
	'command':            '\uE945'
	'compass':            '\uE946'
	'copy':               '\uE947'
	'corner-down-left':   '\uE948'
	'corner-down-right':  '\uE949'
	'corner-left-down':   '\uE94A'
	'corner-left-up':     '\uE94B'
	'corner-right-down':  '\uE94C'
	'corner-right-up':    '\uE94D'
	'corner-up-left':     '\uE94E'
	'corner-up-right':    '\uE94F'
	'cpu':                '\uE950'
	'credit-card':        '\uE951'
	'crop':               '\uE952'
	'crosshair':          '\uE953'
	'database':           '\uE954'
	'delete':             '\uE955'
	'disc':               '\uE956'
	'divide':             '\uE957'
	'divide-circle':      '\uE958'
	'divide-square':      '\uE959'
	'dollar-sign':        '\uE95A'
	'download':           '\uE95B'
	'download-cloud':     '\uE95C'
	'dribbble':           '\uE95D'
	'droplet':            '\uE95E'
	'edit':               '\uE95F'
	'edit-2':             '\uE960'
	'edit-3':             '\uE961'
	'external-link':      '\uE962'
	'eye':                '\uE963'
	'eye-off':            '\uE964'
	'facebook':           '\uE965'
	'fast-forward':       '\uE966'
	'feather':            '\uE967'
	'figma':              '\uE968'
	'file':               '\uE969'
	'file-minus':         '\uE96A'
	'file-plus':          '\uE96B'
	'file-text':          '\uE96C'
	'film':               '\uE96D'
	'filter':             '\uE96E'
	'flag':               '\uE96F'
	'folder':             '\uE970'
	'folder-minus':       '\uE971'
	'folder-plus':        '\uE972'
	'framer':             '\uE973'
	'frown':              '\uE974'
	'gift':               '\uE975'
	'git-branch':         '\uE976'
	'git-commit':         '\uE977'
	'git-merge':          '\uE978'
	'git-pull-request':   '\uE979'
	'github':             '\uE97A'
	'gitlab':             '\uE97B'
	'globe':              '\uE97C'
	'grid':               '\uE97D'
	'hard-drive':         '\uE97E'
	'hash':               '\uE97F'
	'headphones':         '\uE980'
	'heart':              '\uE981'
	'help-circle':        '\uE982'
	'hexagon':            '\uE983'
	'home':               '\uE984'
	'image':              '\uE985'
	'inbox':              '\uE986'
	'info':               '\uE987'
	'instagram':          '\uE988'
	'italic':             '\uE989'
	'key':                '\uE98A'
	'layers':             '\uE98B'
	'layout':             '\uE98C'
	'life-buoy':          '\uE98D'
	'link':               '\uE98E'
	'link-2':             '\uE98F'
	'linkedin':           '\uE990'
	'list':               '\uE991'
	'loader':             '\uE992'
	'lock':               '\uE993'
	'log-in':             '\uE994'
	'log-out':            '\uE995'
	'mail':               '\uE996'
	'map':                '\uE997'
	'map-pin':            '\uE998'
	'maximize':           '\uE999'
	'maximize-2':         '\uE99A'
	'meh':                '\uE99B'
	'menu':               '\uE99C'
	'message-circle':     '\uE99D'
	'message-square':     '\uE99E'
	'mic':                '\uE99F'
	'mic-off':            '\uE9A0'
	'minimize':           '\uE9A1'
	'minimize-2':         '\uE9A2'
	'minus':              '\uE9A3'
	'minus-circle':       '\uE9A4'
	'minus-square':       '\uE9A5'
	'monitor':            '\uE9A6'
	'moon':               '\uE9A7'
	'more-horizontal':    '\uE9A8'
	'more-vertical':      '\uE9A9'
	'mouse-pointer':      '\uE9AA'
	'move':               '\uE9AB'
	'music':              '\uE9AC'
	'navigation':         '\uE9AD'
	'navigation-2':       '\uE9AE'
	'octagon':            '\uE9AF'
	'package':            '\uE9B0'
	'paperclip':          '\uE9B1'
	'pause':              '\uE9B2'
	'pause-circle':       '\uE9B3'
	'pen-tool':           '\uE9B4'
	'percent':            '\uE9B5'
	'phone':              '\uE9B6'
	'phone-call':         '\uE9B7'
	'phone-forwarded':    '\uE9B8'
	'phone-incoming':     '\uE9B9'
	'phone-missed':       '\uE9BA'
	'phone-off':          '\uE9BB'
	'phone-outgoing':     '\uE9BC'
	'pie-chart':          '\uE9BD'
	'play':               '\uE9BE'
	'play-circle':        '\uE9BF'
	'plus':               '\uE9C0'
	'plus-circle':        '\uE9C1'
	'plus-square':        '\uE9C2'
	'pocket':             '\uE9C3'
	'power':              '\uE9C4'
	'printer':            '\uE9C5'
	'radio':              '\uE9C6'
	'refresh-ccw':        '\uE9C7'
	'refresh-cw':         '\uE9C8'
	'repeat':             '\uE9C9'
	'rewind':             '\uE9CA'
	'rotate-ccw':         '\uE9CB'
	'rotate-cw':          '\uE9CC'
	'rss':                '\uE9CD'
	'save':               '\uE9CE'
	'scissors':           '\uE9CF'
	'search':             '\uE9D0'
	'send':               '\uE9D1'
	'server':             '\uE9D2'
	'settings':           '\uE9D3'
	'share':              '\uE9D4'
	'share-2':            '\uE9D5'
	'shield':             '\uE9D6'
	'shield-off':         '\uE9D7'
	'shopping-bag':       '\uE9D8'
	'shopping-cart':      '\uE9D9'
	'shuffle':            '\uE9DA'
	'sidebar':            '\uE9DB'
	'skip-back':          '\uE9DC'
	'skip-forward':       '\uE9DD'
	'slack':              '\uE9DE'
	'slash':              '\uE9DF'
	'sliders':            '\uE9E0'
	'smartphone':         '\uE9E1'
	'smile':              '\uE9E2'
	'speaker':            '\uE9E3'
	'square':             '\uE9E4'
	'star':               '\uE9E5'
	'stop-circle':        '\uE9E6'
	'sun':                '\uE9E7'
	'sunrise':            '\uE9E8'
	'sunset':             '\uE9E9'
	'tablet':             '\uE9EA'
	'tag':                '\uE9EB'
	'target':             '\uE9EC'
	'terminal':           '\uE9ED'
	'thermometer':        '\uE9EE'
	'thumbs-down':        '\uE9EF'
	'thumbs-up':          '\uE9F0'
	'toggle-left':        '\uE9F1'
	'toggle-right':       '\uE9F2'
	'tool':               '\uE9F3'
	'trash':              '\uE9F4'
	'trash-2':            '\uE9F5'
	'trello':             '\uE9F6'
	'trending-down':      '\uE9F7'
	'trending-up':        '\uE9F8'
	'triangle':           '\uE9F9'
	'truck':              '\uE9FA'
	'tv':                 '\uE9FB'
	'twitch':             '\uE9FC'
	'twitter':            '\uE9FD'
	'type':               '\uE9FE'
	'umbrella':           '\uE9FF'
	'underline':          '\uEA00'
	'unlock':             '\uEA01'
	'upload':             '\uEA02'
	'upload-cloud':       '\uEA03'
	'user':               '\uEA04'
	'user-check':         '\uEA05'
	'user-minus':         '\uEA06'
	'user-plus':          '\uEA07'
	'user-x':             '\uEA08'
	'users':              '\uEA09'
	'video':              '\uEA0A'
	'video-off':          '\uEA0B'
	'voicemail':          '\uEA0C'
	'volume':             '\uEA0D'
	'volume-1':           '\uEA0E'
	'volume-2':           '\uEA0F'
	'volume-x':           '\uEA10'
	'watch':              '\uEA11'
	'wifi':               '\uEA12'
	'wifi-off':           '\uEA13'
	'wind':               '\uEA14'
	'x':                  '\uEA15'
	'x-circle':           '\uEA16'
	'x-octagon':          '\uEA17'
	'x-square':           '\uEA18'
	'youtube':            '\uEA19'
	'zap':                '\uEA1A'
	'zap-off':            '\uEA1B'
	'zoom-in':            '\uEA1C'
	'zoom-out':           '\uEA1D'
}
