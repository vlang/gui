module gui

// AlertType configures the type of alert dialog.
//
// - **message** has a title, body and OK button
// - **confirm** is similar to alert but with yes, no buttons
// - **prompt** adds an input field with OK, Cancel buttons
// - **custom** displays the given content. The given content
// is simply displayed. Custom content provides any needed
// callbacks as the standard ones work only for
// the predfined types. See [AlertCfg](#AlertCfg)
pub enum AlertType {
	message
	confirm
	prompt
	custom
}

// AlertCfg configures GUI's alert dialog. [AlertType](#AlertType)
// determines the type of alert. AlertType.message is the default.
// Alerts are asychronous. Keyboard/Mouse input is restricted
// to the alert dialog when visible. Invoke alerts by calling
// [(Window) alert](#Window.alert)
pub struct AlertCfg {
mut:
	visible      bool
	old_id_focus u32
pub:
	alert_type     AlertType
	id             string
	width          f32
	height         f32
	min_width      f32 = 200
	min_height     f32
	max_width      f32 = 300
	max_height     f32
	title          string
	body           string // body text wraps as needed. Newlines supported
	custom_content []View // custom content
	reply          string
	id_focus       u32                     = 7568971
	padding        Padding                 = theme().padding_large
	padding_border Padding                 = theme().padding_border
	on_ok_yes      fn (mut w Window)       = fn (mut _ Window) {}
	on_cancel_no   fn (mut w Window)       = fn (mut _ Window) {}
	on_reply       fn (string, mut Window) = fn (_ string, mut _ Window) {}
}

fn alert_view_generator(cfg AlertCfg) View {
	mut content := []View{}
	content << text(text: cfg.title, text_style: theme().b2)
	content << text(text: cfg.body, wrap: true)
	content << match cfg.alert_type {
		.message { message_view(cfg) }
		.confirm { confirm_view(cfg) }
		.prompt { prompt_view(cfg) }
		.custom { cfg.custom_content }
	}
	return column(
		float:         true
		float_anchor:  .middle_center
		float_tie_off: .middle_center
		color:         theme().color_border
		fill:          true
		padding:       cfg.padding_border
		width:         cfg.width
		height:        cfg.height
		min_width:     cfg.min_width
		max_width:     cfg.max_width
		min_height:    cfg.min_height
		max_height:    cfg.max_height
		content:       [
			column(
				sizing:  fill_fill
				padding: cfg.padding
				h_align: .center
				fill:    true
				color:   theme().color_2
				content: content
			),
		]
	)
}

fn message_view(cfg AlertCfg) []View {
	return [
		button(
			id_focus: cfg.id_focus
			content:  [text(text: 'OK')]
			on_click: fn (_ &ButtonCfg, mut e Event, mut w Window) {
				w.set_id_focus(w.alert_cfg.old_id_focus)
				on_ok_yes := w.alert_cfg.on_ok_yes
				w.alert_cfg = AlertCfg{}
				on_ok_yes(mut w)
				e.is_handled = true
			}
		),
	]
}

fn confirm_view(cfg AlertCfg) []View {
	return [
		row(
			content: [
				button(
					id_focus: cfg.id_focus + 1
					content:  [text(text: 'Yes')]
					on_click: fn (_ &ButtonCfg, mut e Event, mut w Window) {
						w.set_id_focus(w.alert_cfg.old_id_focus)
						on_ok_yes := w.alert_cfg.on_ok_yes
						w.alert_cfg = AlertCfg{}
						on_ok_yes(mut w)
						e.is_handled = true
					}
				),
				button(
					id_focus: cfg.id_focus
					content:  [text(text: 'No')]
					on_click: fn (_ &ButtonCfg, mut e Event, mut w Window) {
						w.set_id_focus(w.alert_cfg.old_id_focus)
						on_cancel_no := w.alert_cfg.on_cancel_no
						w.alert_cfg = AlertCfg{}
						on_cancel_no(mut w)
						e.is_handled = true
					}
				),
			]
		),
	]
}

fn prompt_view(cfg AlertCfg) []View {
	return [
		input(
			id_focus:        cfg.id_focus
			text:            cfg.reply
			sizing:          fill_fit
			on_text_changed: fn (_ &InputCfg, s string, mut w Window) {
				w.alert_cfg = AlertCfg{
					...w.alert_cfg
					reply: s
				}
			}
		),
		row(
			content: [
				button(
					id_focus: cfg.id_focus + 1
					disabled: cfg.reply.len == 0
					content:  [text(text: 'OK')]
					on_click: fn (_ &ButtonCfg, mut e Event, mut w Window) {
						w.set_id_focus(w.alert_cfg.old_id_focus)
						on_reply := w.alert_cfg.on_reply
						reply := w.alert_cfg.reply
						w.alert_cfg = AlertCfg{}
						on_reply(reply, mut w)
						e.is_handled = true
					}
				),
				button(
					id_focus: cfg.id_focus + 2
					content:  [text(text: 'Cancel')]
					on_click: fn (_ &ButtonCfg, mut e Event, mut w Window) {
						w.set_id_focus(w.alert_cfg.old_id_focus)
						on_cancel_no := w.alert_cfg.on_cancel_no
						w.alert_cfg = AlertCfg{}
						on_cancel_no(mut w)
						e.is_handled = true
					}
				),
			]
		),
	]
}
