module markdown

// emoji.v provides emoji shortcode lookup for markdown.
// Supports GitHub-standard shortcodes: :name: -> Unicode emoji.

// emoji_lookup returns the Unicode emoji for a shortcode name,
// or empty string if not found.
pub fn emoji_lookup(name string) string {
	return emoji_map[name] or { '' }
}

// find_emoji_end scans from start for valid emoji shortcode chars.
// Returns end position of name (before closing ':') or -1.
// Max 50 chars scanned. Valid chars: a-z, A-Z, 0-9, _, +, -.
// First char must be alpha, underscore, + or -.
pub fn find_emoji_end(text string, start int) int {
	if start >= text.len {
		return -1
	}
	// First char: alpha, underscore, + or -
	fc := text[start]
	if !((fc >= `a` && fc <= `z`) || (fc >= `A` && fc <= `Z`) || fc == `_` || fc == `+` || fc == `-`) {
		return -1
	}
	mut i := start + 1
	limit := if start + 50 < text.len { start + 50 } else { text.len }
	for i < limit {
		ch := text[i]
		if ch == `:` {
			return i
		}
		if (ch >= `a` && ch <= `z`) || (ch >= `A` && ch <= `Z`)
			|| (ch >= `0` && ch <= `9`) || ch == `_` || ch == `+` || ch == `-` {
			i++
			continue
		}
		return -1 // invalid char
	}
	return -1
}

// emoji_map maps GitHub-standard shortcode names to Unicode emoji.
const emoji_map = {
	// Smileys & Emotion
	'smile':                        '😄'
	'laughing':                     '😆'
	'blush':                        '😊'
	'smiley':                       '😃'
	'grinning':                     '😀'
	'grin':                         '😁'
	'joy':                          '😂'
	'rofl':                         '🤣'
	'sweat_smile':                  '😅'
	'wink':                         '😉'
	'kissing_heart':                '😘'
	'yum':                          '😋'
	'stuck_out_tongue':             '😛'
	'stuck_out_tongue_winking_eye': '😜'
	'stuck_out_tongue_closed_eyes': '😝'
	'sunglasses':                   '😎'
	'heart_eyes':                   '😍'
	'thinking':                     '🤔'
	'neutral_face':                 '😐'
	'expressionless':               '😑'
	'unamused':                     '😒'
	'sweat':                        '😓'
	'pensive':                      '😔'
	'confused':                     '😕'
	'confounded':                   '😖'
	'disappointed':                 '😞'
	'worried':                      '😟'
	'angry':                        '😠'
	'rage':                         '😡'
	'cry':                          '😢'
	'sob':                          '😭'
	'fearful':                      '😨'
	'scream':                       '😱'
	'tired_face':                   '😫'
	'sleeping':                     '😴'
	'sleepy':                       '😪'
	'mask':                         '😷'
	'nerd_face':                    '🤓'
	'cowboy_hat_face':              '🤠'
	'clown_face':                   '🤡'
	'nauseated_face':               '🤢'
	'rolling_eyes':                 '🙄'
	'hushed':                       '😯'
	'frowning':                     '😦'
	'anguished':                    '😧'
	'imp':                          '👿'
	'smiling_imp':                  '😈'
	'skull':                        '💀'
	'ghost':                        '👻'
	'alien':                        '👾'
	'robot':                        '🤖'
	'poop':                         '💩'
	'hankey':                       '💩'
	'clap':                         '👏'
	'wave':                         '👋'
	'raised_hands':                 '🙌'
	'pray':                         '🙏'
	'handshake':                    '🤝'
	'muscle':                       '💪'
	'point_up':                     '☝️'
	'point_down':                   '👇'
	'point_left':                   '👈'
	'point_right':                  '👉'
	'middle_finger':                '🖕'
	'raised_hand':                  '✋'
	'ok_hand':                      '👌'
	'thumbsup':                     '👍'
	'thumbsdown':                   '👎'
	'fist':                         '✊'
	'punch':                        '👊'
	'v':                            '✌️'
	'crossed_fingers':              '🤞'
	'metal':                        '🤘'
	'eyes':                         '👀'
	'tongue':                       '👅'
	'lips':                         '👄'
	// Hearts & Symbols
	'heart':                        '❤️'
	'yellow_heart':                 '💛'
	'green_heart':                  '💚'
	'blue_heart':                   '💙'
	'purple_heart':                 '💜'
	'black_heart':                  '🖤'
	'broken_heart':                 '💔'
	'heartbeat':                    '💓'
	'heartpulse':                   '💗'
	'sparkling_heart':              '💖'
	'cupid':                        '💘'
	'gift_heart':                   '💝'
	'heart_decoration':             '💟'
	'sparkles':                     '✨'
	'star':                         '⭐'
	'star2':                        '🌟'
	'dizzy':                        '💫'
	'boom':                         '💥'
	'fire':                         '🔥'
	'droplet':                      '💧'
	'100':                          '💯'
	'zap':                          '⚡'
	'snowflake':                    '❄️'
	'rainbow':                      '🌈'
	'sun_with_face':                '🌞'
	'cloud':                        '☁️'
	'umbrella':                     '☂️'
	// People
	'baby':                         '👶'
	'boy':                          '👦'
	'girl':                         '👧'
	'man':                          '👨'
	'woman':                        '👩'
	'older_man':                    '👴'
	'older_woman':                  '👵'
	// Animals
	'dog':                          '🐶'
	'cat':                          '🐱'
	'mouse':                        '🐭'
	'hamster':                      '🐹'
	'rabbit':                       '🐰'
	'fox_face':                     '🦊'
	'bear':                         '🐻'
	'panda_face':                   '🐼'
	'koala':                        '🐨'
	'tiger':                        '🐯'
	'lion':                         '🦁'
	'cow':                          '🐮'
	'pig':                          '🐷'
	'frog':                         '🐸'
	'monkey_face':                  '🐵'
	'see_no_evil':                  '🙈'
	'hear_no_evil':                 '🙉'
	'speak_no_evil':                '🙊'
	'chicken':                      '🐔'
	'penguin':                      '🐧'
	'bird':                         '🐦'
	'eagle':                        '🦅'
	'butterfly':                    '🦋'
	'bug':                          '🐛'
	'snail':                        '🐌'
	'snake':                        '🐍'
	'turtle':                       '🐢'
	'octopus':                      '🐙'
	'whale':                        '🐳'
	'dolphin':                      '🐬'
	'fish':                         '🐟'
	'unicorn':                      '🦄'
	'bee':                          '🐝'
	'crab':                         '🦀'
	// Food & Drink
	'apple':                        '🍎'
	'green_apple':                  '🍏'
	'banana':                       '🍌'
	'grapes':                       '🍇'
	'watermelon':                   '🍉'
	'strawberry':                   '🍓'
	'peach':                        '🍑'
	'cherries':                     '🍒'
	'pineapple':                    '🍍'
	'lemon':                        '🍋'
	'avocado':                      '🥑'
	'pizza':                        '🍕'
	'hamburger':                    '🍔'
	'fries':                        '🍟'
	'hotdog':                       '🌭'
	'taco':                         '🌮'
	'burrito':                      '🌯'
	'egg':                          '🥚'
	'coffee':                       '☕'
	'tea':                          '🍵'
	'beer':                         '🍺'
	'wine_glass':                   '🍷'
	'cocktail':                     '🍸'
	'cake':                         '🍰'
	'cookie':                       '🍪'
	'chocolate_bar':                '🍫'
	'candy':                        '🍬'
	'ice_cream':                    '🍨'
	'doughnut':                     '🍩'
	// Objects
	'computer':                     '💻'
	'keyboard':                     '⌨️'
	'phone':                        '☎️'
	'iphone':                       '📱'
	'envelope':                     '✉️'
	'email':                        '📧'
	'inbox_tray':                   '📥'
	'outbox_tray':                  '📤'
	'package':                      '📦'
	'memo':                         '📝'
	'pencil2':                      '✏️'
	'book':                         '📖'
	'books':                        '📚'
	'bookmark':                     '🔖'
	'link':                         '🔗'
	'paperclip':                    '📎'
	'scissors':                     '✂️'
	'lock':                         '🔒'
	'unlock':                       '🔓'
	'key':                          '🔑'
	'hammer':                       '🔨'
	'wrench':                       '🔧'
	'gear':                         '⚙️'
	'bulb':                         '💡'
	'flashlight':                   '🔦'
	'battery':                      '🔋'
	'mag':                          '🔍'
	'mag_right':                    '🔎'
	'bell':                         '🔔'
	'no_bell':                      '🔕'
	'loudspeaker':                  '📢'
	'mega':                         '📣'
	'mute':                         '🔇'
	'speaker':                      '🔈'
	'sound':                        '🔉'
	'loud_sound':                   '🔊'
	'hourglass':                    '⌛'
	'alarm_clock':                  '⏰'
	'watch':                        '⌚'
	'calendar':                     '📅'
	'chart':                        '📈'
	'chart_with_downwards_trend':   '📉'
	'bar_chart':                    '📊'
	'clipboard':                    '📋'
	'pushpin':                      '📌'
	'round_pushpin':                '📍'
	'triangular_flag_on_post':      '🚩'
	'trophy':                       '🏆'
	'medal_sports':                 '🏅'
	'1st_place_medal':              '🥇'
	'2nd_place_medal':              '🥈'
	'3rd_place_medal':              '🥉'
	'crown':                        '👑'
	'gem':                          '💎'
	'moneybag':                     '💰'
	'dollar':                       '💵'
	'credit_card':                  '💳'
	'gift':                         '🎁'
	'balloon':                      '🎈'
	'tada':                         '🎉'
	'confetti_ball':                '🎊'
	'rocket':                       '🚀'
	'airplane':                     '✈️'
	'car':                          '🚗'
	'bus':                          '🚌'
	'train':                        '🚆'
	'bike':                         '🚲'
	'ship':                         '🚢'
	'anchor':                       '⚓'
	'earth_americas':               '🌎'
	'earth_africa':                 '🌍'
	'earth_asia':                   '🌏'
	'globe_with_meridians':         '🌐'
	'house':                        '🏠'
	'office':                       '🏢'
	'hospital':                     '🏥'
	'school':                       '🏫'
	// Symbols & Signs
	'white_check_mark':             '✅'
	'ballot_box_with_check':        '☑️'
	'heavy_check_mark':             '✔️'
	'x':                            '❌'
	'negative_squared_cross_mark':  '❎'
	'bangbang':                     '‼️'
	'interrobang':                  '⁉️'
	'question':                     '❓'
	'grey_question':                '❔'
	'grey_exclamation':             '❕'
	'exclamation':                  '❗'
	'warning':                      '⚠️'
	'no_entry':                     '⛔'
	'no_entry_sign':                '🚫'
	'stop_sign':                    '🛑'
	'construction':                 '🚧'
	'recycle':                      '♻️'
	'information_source':           'ℹ️'
	'sos':                          '🆘'
	'new':                          '🆕'
	'up':                           '🆙'
	'cool':                         '🆒'
	'free':                         '🆓'
	'ok':                           '🆗'
	'arrow_up':                     '⬆️'
	'arrow_down':                   '⬇️'
	'arrow_left':                   '⬅️'
	'arrow_right':                  '➡️'
	'arrow_upper_right':            '↗️'
	'arrow_lower_right':            '↘️'
	'arrow_lower_left':             '↙️'
	'arrow_upper_left':             '↖️'
	'arrows_counterclockwise':      '🔄'
	'leftwards_arrow_with_hook':    '↩️'
	'arrow_right_hook':             '↪️'
	'ten':                          '🔟'
	'copyright':                    '©️'
	'registered':                   '®️'
	'tm':                           '™️'
	// Flags (common)
	'checkered_flag':               '🏁'
	'white_flag':                   '🏳️'
	// Common aliases
	'+1':                           '👍'
	'-1':                           '👎'
}
