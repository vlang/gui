module gui

// AI-DOC: window_update.v
// - Scope: Window frame/update/render pipeline.
// - Entry points: frame_fn() from gg, update_view(), update_window().
// - Refresh flags: layout refresh overrides render-only refresh.
// - Order: init subsystems -> flush commands -> update/layout/renderers ->
//   run SVG offscreen filter passes -> draw swapchain pass.
// - Locking: layout/renderer rebuild runs under window lock.
import log
import sokol.sapp

// frame_fn is the only place where the window is rendered.
// see: CLAUDE.md §Render Pipeline for the full flow diagram.
fn frame_fn(mut window Window) {
	window.init_ime()
	window.init_a11y()
	window.flush_commands()

	if window.refresh_layout {
		window.update()
		window.sync_a11y()
		window.refresh_layout = false
		window.refresh_render_only = false
	} else if window.refresh_render_only {
		window.update_render_only()
		window.refresh_render_only = false
	}

	// Process SVG filters in offscreen passes BEFORE the
	// swapchain pass; sokol doesn't support nested passes.
	process_svg_filters(mut window)

	window.lock()
	window.ui.begin()
	renderers_draw(mut window)
	window.ui.end()
	window.unlock()
	sapp.set_mouse_cursor(window.view_state.mouse_cursor)
}

// update_view replaces the current view generator and clears view state.
pub fn (mut window Window) update_view(gen_view fn (&Window) View) {
	window.lock()
	window.clear_view_state()
	window.view_generator = gen_view
	window.unlock()
	window.update_window()
}

// update_window marks the window as needing an update. The actual update
// (re-calculating layout and generating renderers) is performed at the start
// of the next frame to batch multiple state changes.
pub fn (mut window Window) update_window() {
	window.mark_layout_refresh()
	window.ui.refresh_ui()
}

fn (mut window Window) request_render_only() {
	window.mark_render_only_refresh()
	window.ui.refresh_ui()
}

fn (mut window Window) mark_layout_refresh() {
	window.refresh_layout = true
	window.refresh_render_only = false
}

fn (mut window Window) mark_render_only_refresh() {
	if !window.refresh_layout {
		window.refresh_render_only = true
	}
}

// update generates a new layout from the window's current view generator.
fn (mut window Window) update() {
	log.debug('update_window')
	//--------------------------------------------
	window.lock()
	clip_rect := window.window_rect()
	background_color := window.color_background()

	mut view := window.view_generator(window)
	$if !prod {
		if window.inspector_enabled {
			window.inspector_props_cache = map[string]InspectorNodeProps{}
			selected := inspector_selected_path(window)
			window.inspector_tree_cache = inspector_build_tree_nodes(&window.layout, selected, mut
				window.inspector_props_cache)
		}
	}
	layout_clear(mut window.layout)
	window.layout = window.compose_layout(mut view)
	window.build_renderers(background_color, clip_rect)
	window.unlock()
	//--------------------------------------------

	view_clear(mut view)
	window.stats.update_max_renderers(usize(window.renderers.len))
}

fn (mut window Window) update_render_only() {
	log.debug('update_render_only')
	//--------------------------------------------
	window.lock()
	clip_rect := window.window_rect()
	background_color := window.color_background()
	window.build_renderers(background_color, clip_rect)
	window.unlock()
	//--------------------------------------------

	window.stats.update_max_renderers(usize(window.renderers.len))
}

fn (mut window Window) build_renderers(background_color Color, clip_rect DrawClip) {
	// process_svg_filters swaps renderer buffers. Reset both
	// arrays before render so buffers are reused safely.
	mut filter_renderers := window.scratch.take_filter_renderers(0)
	window.scratch.put_filter_renderers(mut filter_renderers)
	window.scratch.begin_svg_transform_batches()
	array_clear(mut window.renderers)
	render_layout(mut window.layout, background_color, clip_rect, mut window)
	window.scratch.trim_svg_transform_batches()
	$if !prod {
		if window.inspector_enabled {
			inspector_inject_wireframe(mut window)
		}
	}

	// Render RTF tooltip if active
	if window.view_state.rtf_tooltip_text != '' {
		window.render_rtf_tooltip(clip_rect)
	}
}

// compose_layout takes the View generated by the user's view function and
// processes it into a fully resolved Layout tree. This involves:
// 1. Transforming the View tree into a Layout tree (`generate_layout`)
// 2. Calculating sizes and positions for all elements (`layout_arrange`)
// 3. Wrapping the result in a root Layout with a transparent background
fn (mut window Window) compose_layout(mut view View) Layout {
	timer := if window.debug_layout { layout_stats_timer_start() } else { LayoutStatsTimer{} }

	mut layout := generate_layout(mut view, mut window)
	// amend_layout callbacks fire inside layout_arrange (during size/position
	// passes), NOT during render_layout. See CLAUDE.md §Layout Pipeline.
	layouts := layout_arrange(mut layout, mut window)
	result := Layout{
		shape:    &Shape{
			color: color_transparent
		}
		children: layouts
	}

	if window.debug_layout {
		window.layout_stats = LayoutStats{
			total_time_us:  timer.elapsed_us()
			node_count:     count_nodes(&result)
			floating_count: layouts.len - 1
		}
	}

	return result
}
