module gui

pub struct TextSpan {
	id    string
	text  string
	style TextStyle
	x     f32
	y     f32
}
