module titlebar

pub fn prefer_dark_titlebar(handle voidptr, dark bool) {}
